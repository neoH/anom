/*
This module can be divided into several sub modules: issue module, computing module and retiring module.
*/
module ieu (
	);






endmodule
