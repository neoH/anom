/*********************************************************************************************
*********************************************************************************************/
module anom(

);


// instantiating sub modules of anom

// interface module, which used to translate self-defined communication protocol to public
// interface protocols.



endmodule
