/*
This module can be divided into several sub modules: issue module, computing module and retiring module.
----------------------------------------------------------------------------------------------------------
Interface Protocol:
----------------------------------------------------------------------------------------------------------
*/
module ieu (
	);






endmodule
