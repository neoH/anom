/*
The assertion block for ifu module
*/

module ifu_ast_block(
	input logic i_Clk,
);



endmodule
