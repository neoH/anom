module ieu (
	);


endmodule
